class common;

  static mailbox gen2drv = new();
  static virtual sp_intf intf;
  static mailbox mon2scb = new();

endclass
